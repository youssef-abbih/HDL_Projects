library verilog;
use verilog.vl_types.all;
entity multiplication_vlg_vec_tst is
end multiplication_vlg_vec_tst;
